parameter off          = 7'b1111111;

parameter PLL_Locked   = 7'b1000111;
parameter PLL_Unlocked = 7'b1000001;

parameter top          = 7'b1111110;
parameter upper_right  = 7'b1111101;
parameter lower_right  = 7'b1111011;
parameter bottom       = 7'b1110111;

