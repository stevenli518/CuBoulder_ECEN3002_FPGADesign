`ifndef _parameter_vh_
`define _parameter_vh_
//Horizontal Parameters
parameter Total_Pixels = 800;
parameter Active_Pixel =640;
parameter H_Front_P =16;
parameter H_Back_P=48;
parameter H_Sync_W = 96;

//Vertical Parameters
parameter Total_lines = 525;
parameter Active_Line = 480;
parameter V_Front_P =10;
parameter V_Back_P=33;
parameter V_Sync_W = 2;
`endif