`ifndef _parameter_vh_
`define _parameter_vh_
//Horizontal Parameters
parameter Total_Pixels = 1650;
parameter Active_Pixel =1280;
parameter H_Front_P =110;
parameter H_Back_P=220;
parameter H_Sync_W = 40;

//Vertical Parameters
parameter Total_lines = 750;
parameter Active_Line = 720;
parameter V_Front_P =5;
parameter V_Back_P=20;
parameter V_Sync_W = 5;
`endif